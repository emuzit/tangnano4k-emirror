//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07 Education
//Part Number: GW1NSR-LV4CQN48PC6/I5
//Device: GW1NSR-4C
//Created Time: Fri Oct 28 12:25:59 2022

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [8:0] ad;

wire [15:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[15:0],dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({gw_gnd,ad[8:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "ASYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0018303400FF301800FF30170020474000033103004230080082300800113103;
defparam prom_inst_0.INIT_RAM_01 = 256'h00A0370400E036210012363300E23632000E3631003636300001310800043037;
defparam prom_inst_0.INIT_RAM_02 = 256'h000A39010010390600023905001A37050060370B0001371700783715005A3703;
defparam prom_inst_0.INIT_RAM_03 = 256'h00433A130050471C0020371B005236200060302D003336010008360000123731;
defparam prom_inst_0.INIT_RAM_04 = 256'h00283C0400343C010001362200403634000336360013363500F83A1900003A18;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000381000403C0B009C3C0A001C3C0900003C0800083C0700003C0600983C05;
defparam prom_inst_0.INIT_RAM_06 = 256'h0058300E00FF300400003000001A400500024001006437080000381200103811;
defparam prom_inst_0.INIT_RAM_07 = 256'h00303A1B00283A1000303A0F00A750000000440E0001501F006143000000302E;
defparam prom_inst_0.INIT_RAM_08 = 256'h00125804000F5803000F5802001458010023580000143A1F00603A1100263A1E;
defparam prom_inst_0.INIT_RAM_09 = 256'h0008580C000D580B0008580A000558090005580800085807000C580600265805;
defparam prom_inst_0.INIT_RAM_0A = 256'h00005814000358130007581200095811000358100000580F0000580E0003580D;
defparam prom_inst_0.INIT_RAM_0B = 256'h0008581C0006581B0005581A00085819000D5818000858170003581600015815;
defparam prom_inst_0.INIT_RAM_0C = 256'h00465824002858230015582200115821001158200017581F0029581E000E581D;
defparam prom_inst_0.INIT_RAM_0D = 256'h0024582C0022582B0024582A0026582900645828002658270008582600265825;
defparam prom_inst_0.INIT_RAM_0E = 256'h00245834002658330024583200425831004058300022582F0006582E0024582D;
defparam prom_inst_0.INIT_RAM_0F = 256'h0042583C0028583B0026583A0024583900445838002658370022583600225835;
defparam prom_inst_0.INIT_RAM_10 = 256'h000951860024518500255184001451830000518200F2518100FF518000CE583D;
defparam prom_inst_0.INIT_RAM_11 = 256'h003D518E0042518D00B2518C00E0518B0054518A007551890009518800095187;
defparam prom_inst_0.INIT_RAM_12 = 256'h0003519600F0519500F05194007051930004519200F85191004651900056518F;
defparam prom_inst_0.INIT_RAM_13 = 256'h0038519E0082519D0006519C0000519B0004519A001251990004519800015197;
defparam prom_inst_0.INIT_RAM_14 = 256'h007D548700715486006554850051548400285483001454820008548100015480;
defparam prom_inst_0.INIT_RAM_15 = 256'h00EA548F00DD548E00CD548D00B8548C00AA548B009A548A0091548900875488;
defparam prom_inst_0.INIT_RAM_16 = 256'h007C538700885386007E5385000A538400085383005B5382001E5381001D5490;
defparam prom_inst_0.INIT_RAM_17 = 256'h001055890010558400405583000655800098538B0001538A00105389006C5388;
defparam prom_inst_0.INIT_RAM_18 = 256'h00085304000053030010530200305301000853000040501D00F8558B0000558A;
defparam prom_inst_0.INIT_RAM_19 = 256'h000050250006530C0004530B0030530A00085309001653070008530600305305;
defparam prom_inst_0.INIT_RAM_1A = 256'h0031381500313814000738210047382000073C07006330360011303500023008;
defparam prom_inst_0.INIT_RAM_1B = 256'h00A9380700063806003F3805000A380400FA3803000038020000380100003800;
defparam prom_inst_0.INIT_RAM_1C = 256'h00EE380F0002380E0072380D0006380C00D0380B0002380A0000380900053808;
defparam prom_inst_0.INIT_RAM_1D = 256'h00E03A1500023A1400023A020003370C00523709002936120000361800043813;
defparam prom_inst_0.INIT_RAM_1E = 256'h001648370020460C0037460B000444070003471300C33006001C300200024004;
defparam prom_inst_0.INIT_RAM_1F = 256'h00000000000000000000000000000000FFFFFFFF000035030083500100043824;

endmodule //Gowin_pROM
